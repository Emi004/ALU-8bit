module alu (
);
    
endmodule