`include "cu.v"
`include "au.v"

module alu (
    input clk,rst,
    input [1:0] select,
    input [7:0]A,B,
    output[15:0] result,
    output overflow,negative,zero,carry_out,divisionBy0,done
);
    
    wire startadd,startsub,startmultiplier,startdiv;
    cu CU(.done(done),.clk(clk),.rst(rst),.s(select),.startadd(startadd),.startsub(startsub),.startdiv(startdiv),.startmultiplier(startmultiplier));
    au AU(.clk(clk),.rst(rst),.A(A),.B(B),.startadd(startadd),.startsub(startsub),
        .startdiv(startdiv),.startmultiplier(startmultiplier),.result(result),
        .overflow(overflow),.negative(negative),.zero(zero),.carry_out(carry_out),.divisionBy0(divisionBy0),
        .done(done)
    );

endmodule

`timescale 1ns/1ps

module alu_tb;

    // Inputs
    reg clk;
    reg rst;
    reg [1:0] select;
    reg [7:0] A;
    reg [7:0] B;

    // Outputs
    wire [15:0] result;
    wire overflow, negative, zero, carry_out, divisionBy0, done;

    // Instantiate the ALU
    alu uut (
        .clk(clk),
        .rst(rst),
        .select(select),
        .A(A),
        .B(B),
        .result(result),
        .overflow(overflow),
        .negative(negative),
        .zero(zero),
        .carry_out(carry_out),
        .divisionBy0(divisionBy0),
        .done(done)
    );

    // Clock generation (100MHz)
    initial begin
        clk = 0;
        rst = 1;
        
        #10 rst = 0; // Release reset after 5 time units
        forever #5 clk = ~clk;
    end
    initial begin
    // Wait after reset
    #10;

    // Addition test
    select = 2'b00; A = 8'd15; B = 8'd8;
    wait(done); @(posedge clk); wait(!done);
    $display("Addition:       A = %0d, B = %0d, Result = %0d, Overflow = %b, Negative = %b, Zero = %b, Carry Out = %b", A, B, result[7:0], overflow, negative, zero, carry_out);

    // Subtraction test
    select = 2'b01; A = 8'd15; B = 8'd8;
    wait(done); @(posedge clk); wait(!done);
    $display("Subtraction:    A = %0d, B = %0d, Result = %0d, Overflow = %b, Negative = %b, Zero = %b, Carry Out = %b", A, B, result[7:0], overflow, negative, zero, carry_out);

    // Multiplication test
    select = 2'b10; A = 8'd15; B = 8'd8;
    wait(done); @(posedge clk); wait(!done);
    $display("Multiplication: A = %0d, B = %0d, Result = %0d, Overflow = %b, Negative = %b, Zero = %b, Carry Out = %b", A, B, result, overflow, negative, zero, carry_out);

    // Division test
    select = 2'b11; A = 8'd15; B = 8'd8;
    wait(done); @(posedge clk); wait(!done);
    $display("Division:       A = %0d, B = %0d, Result = %0d, Reminder=%0d, Overflow = %b, Negative = %b, Zero = %b, Carry Out = %b,div 0 = %b", A, B, result[15:8], result[7:0],overflow, negative, zero, carry_out,divisionBy0);

    // Division 0 test
    select = 2'b11; A = 8'd15; B = 8'd0;
    wait(done); @(posedge clk); wait(!done);
    $display("Division:       A = %0d, B = %0d, Result = %0d, Reminder=%0d, Overflow = %b, Negative = %b, Zero = %b, Carry Out = %b,div 0=%b", A, B, result[15:8], result[7:0],overflow, negative, zero, carry_out, divisionBy0);

    $finish;
end

         

endmodule
